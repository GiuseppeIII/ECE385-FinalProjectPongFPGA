//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 298 Lab 7                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball ( input Reset, frame_clk,
					input [7:0] keycode,
					input	[9:0] Paddle1X, Paddle1Y, Paddle2X, Paddle2Y, 
									Paddle1L, Paddle1W, Paddle2L, Paddle2W,	
               output [9:0]  BallX, BallY, BallS );
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion, Ball_Size;
	 
    parameter [9:0] Ball_X_Center=320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center=240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min=33;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max=596;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min=20;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max=461;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step=4;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step=4;      // Step size on the Y axis

    assign Ball_Size = 4;  // assigns the value 4 as a 10-digit binary number, ie "0000000100"
	 int paddle1minHeight, paddle1maxHeight, paddle1minWidth, paddle1maxWidth;
	 int paddle2minHeight, paddle2maxHeight, paddle2minWidth, paddle2maxWidth;
	 int ballymotion, bally2motion;
	 
	 assign paddle1minHeight = Paddle1Y - Paddle1L;
	 assign paddle1maxHeight = Paddle1Y + Paddle1L;
	 assign paddle1minWidth = Paddle1X - Paddle1W;
	 assign paddle1maxWidth = Paddle1X + Paddle1W;
	 
	 assign paddle2minHeight = Paddle2Y - Paddle2L;
	 assign paddle2maxHeight = Paddle2Y + Paddle2L;
	 assign paddle2minWidth = Paddle2X - Paddle2W;
	 assign paddle2maxWidth = Paddle2X + Paddle2W;
	 
	 assign bally1motion = (Ball_Y_Pos - Paddle1Y)>>3;
	 assign bally2motion = (Ball_Y_Pos - Paddle2Y)>>3;
   
    always_ff @ (posedge Reset or posedge frame_clk )
    begin: Move_Ball
        if (Reset)  // Asynchronous Reset
		  //initalize ball
        begin 
            Ball_Y_Motion <= 0;
				Ball_X_Motion <= Ball_X_Step;
				Ball_Y_Pos <= Ball_Y_Center;
				Ball_X_Pos <= Ball_X_Center;
        end
           
        else 
        begin 
				Ball_Y_Motion <= Ball_Y_Motion;
				
				if ( (Ball_Y_Pos + Ball_Size) >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
					  Ball_Y_Motion <= (~ (Ball_Y_Step) + 1'b1);  // 2's complement. 
				 
				else if ( (Ball_Y_Pos - Ball_Size) <= Ball_Y_Min )  // Ball is at the top edge, BOUNCE!
					  Ball_Y_Motion <= Ball_Y_Step;
					    
				else if ( (Ball_X_Pos + Ball_Size) >= Ball_X_Max )  // Ball is at the Right edge, BOUNCE!
					  Ball_X_Motion <= (~ (Ball_X_Step) + 1'b1);  // 2's complement.
					  	  
				else if ( (Ball_X_Pos - Ball_Size) <= Ball_X_Min )  // Ball is at the Left edge, BOUNCE!
					  Ball_X_Motion <= Ball_X_Step;
					 
				//if hits paddle1
				//rightEdge
				if (((Ball_X_Pos - Ball_Size) <= paddle1maxWidth) && 
					((Ball_Y_Pos - Ball_Size) <= paddle1maxHeight ) &&
					((Ball_Y_Pos + Ball_Size) >= paddle1minHeight ))
					begin
						Ball_X_Motion <= Ball_X_Step;
						Ball_Y_Motion <= bally1motion;
						if (bally1motion < 0)
							Ball_Y_Motion <= (~ (bally1motion) + 1'b1);
					end
				
				//if hits paddle2
				//leftEdge
				if (((Ball_X_Pos + Ball_Size) >= paddle2minWidth) && 
					((Ball_Y_Pos - Ball_Size) <= paddle2maxHeight ) &&
					((Ball_Y_Pos + Ball_Size) >= paddle2minHeight ))
					begin
						Ball_X_Motion <= (~ (Ball_X_Step) + 1'b1);
						Ball_Y_Motion <= bally2motion;
						if (bally2motion < 0)
							Ball_Y_Motion <= (~ (bally2motion) + 1'b1);
					end
				
//				 case (keycode)
//					8'h04 : begin
//								if ((Ball_X_Pos - Ball_Size) > Ball_X_Min)
//									begin
//										Ball_X_Motion <= -Ball_X_Step;//A
//										Ball_Y_Motion<= 0;
//									end
//							  end    
//					8'h07 : begin
//								if ((Ball_X_Pos + Ball_Size) < Ball_X_Max)
//									begin	
//										Ball_X_Motion <= Ball_X_Step;//D
//										Ball_Y_Motion <= 0;	
//									end
//							  end 
//					8'h16 : begin
//								if ((Ball_Y_Pos + Ball_Size) < Ball_Y_Max)
//									begin	
//										Ball_Y_Motion <= Ball_Y_Step;//S
//										Ball_X_Motion <= 0;		
//									end   
//							 end		  
//					8'h1A : begin
//								if ((Ball_Y_Pos - Ball_Size) > Ball_Y_Min)
//									begin
//										Ball_Y_Motion <= -Ball_Y_Step;//W
//										Ball_X_Motion <= 0;
//									end
//							 end	  
//					default: ;
//			   endcase
				 
				Ball_Y_Pos <= (Ball_Y_Pos + Ball_Y_Motion);  // Update ball position
				Ball_X_Pos <= (Ball_X_Pos + Ball_X_Motion);
			
		end  
    end
       
    assign BallX = Ball_X_Pos;
    assign BallY = Ball_Y_Pos;
    assign BallS = Ball_Size;

endmodule
