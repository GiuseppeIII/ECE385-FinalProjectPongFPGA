module font_rom ( input [8:0]	addr,
						output [31:0]	data
					 );

	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
			// code x00
        32'b00000000000000000000000000000000, // 00 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 01 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 02 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 03 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 04 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 05 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 06 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 07 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 08 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 09 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 0a ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 0b ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 0c ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 0d ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 0e ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 0f ||||||||||||||||||||||||||||||||
		  32'b11111111000000000000111111110000, // 10 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 11 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 12 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 13 ||||||||||||||||||||||||||||||||
        32'b11111111000000001111111111110000, // 14 ||||||||||||||||||||||||||||||||
        32'b11111111000000001111111111110000, // 15 ||||||||||||||||||||||||||||||||
        32'b11111111000000001111111111110000, // 16 ||||||||||||||||||||||||||||||||
        32'b11111111000000001111111111110000, // 17 ||||||||||||||||||||||||||||||||
        32'b11111111000011111111111111110000, // 18 ||||||||||||||||||||||||||||||||
        32'b11111111000011111111111111110000, // 19 ||||||||||||||||||||||||||||||||
        32'b11111111000011111111111111110000, // 1a ||||||||||||||||||||||||||||||||
        32'b11111111000011111111111111110000, // 1b ||||||||||||||||||||||||||||||||
        32'b11111111111111110000111111110000, // 1c ||||||||||||||||||||||||||||||||
        32'b11111111111111110000111111110000, // 1d ||||||||||||||||||||||||||||||||
        32'b11111111111111110000111111110000, // 1e ||||||||||||||||||||||||||||||||
        32'b11111111111111110000111111110000, // 1f ||||||||||||||||||||||||||||||||
		  32'b11111111111100000000111111110000, // 20 ||||||||||||||||||||||||||||||||
        32'b11111111111100000000111111110000, // 21 ||||||||||||||||||||||||||||||||
        32'b11111111111100000000111111110000, // 22 ||||||||||||||||||||||||||||||||
        32'b11111111111100000000111111110000, // 23 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 24 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 25 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 26 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 27 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 28 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 29 ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 2a ||||||||||||||||||||||||||||||||
        32'b11111111000000000000111111110000, // 2b ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 2c ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 2d ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 2e ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111100000000, // 2f ||||||||||||||||||||||||||||||||
		  32'b00000000000000000000000000000000, // 30 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 31 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 32 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 33 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 34 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 35 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 36 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 37 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 38 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 39 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3a ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3b ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3c ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3d ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3e ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3f |||||||||||||||||||||||||||||||| 
         // code x01
        32'b00000000000000000000000000000000, // 00 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 01 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 02 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 03 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 04 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 05 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 06 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 07 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 08 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 09 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 0a ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 0b ||||||||||||||||||||||||||||||||
        32'b00000000111111111111000000000000, // 0c ||||||||||||||||||||||||||||||||
        32'b00000000111111111111000000000000, // 0d ||||||||||||||||||||||||||||||||
        32'b00000000111111111111000000000000, // 0e ||||||||||||||||||||||||||||||||
        32'b00000000111111111111000000000000, // 0f ||||||||||||||||||||||||||||||||
		  32'b00001111111111111111000000000000, // 10 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111000000000000, // 11 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111000000000000, // 12 ||||||||||||||||||||||||||||||||
        32'b00001111111111111111000000000000, // 13 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 14 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 15 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 16 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 17 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 18 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 19 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1a ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1b ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1c ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1d ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1e ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 1f ||||||||||||||||||||||||||||||||
		  32'b00000000000011111111000000000000, // 20 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 21 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 22 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 23 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 24 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 25 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 26 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 27 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 28 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 29 ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 2a ||||||||||||||||||||||||||||||||
        32'b00000000000011111111000000000000, // 2b ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111111110000, // 2c ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111111110000, // 2d ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111111110000, // 2e ||||||||||||||||||||||||||||||||
        32'b00001111111111111111111111110000, // 2f ||||||||||||||||||||||||||||||||
		  32'b00000000000000000000000000000000, // 30 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 31 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 32 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 33 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 34 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 35 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 36 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 37 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 38 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 39 ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3a ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3b ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3c ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3d ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3e ||||||||||||||||||||||||||||||||
        32'b00000000000000000000000000000000, // 3f ||||||||||||||||||||||||||||||||
         // code x02
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
         // code x03
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
         // code x04
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000011111111111100000000,
32'b00000000000011111111111100000000,
32'b00000000000011111111111100000000,
32'b00000000000011111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00000000111111111111111100000000,
32'b00001111111100001111111100000000,
32'b00001111111100001111111100000000,
32'b00001111111100001111111100000000,
32'b00001111111100001111111100000000,
32'b11111111000000001111111100000000,
32'b11111111000000001111111100000000,
32'b11111111000000001111111100000000,
32'b11111111000000001111111100000000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000011111111111111110000,
32'b00000000000011111111111111110000,
32'b00000000000011111111111111110000,
32'b00000000000011111111111111110000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
         // code x05
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
         // code x06
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000111111111111000000000000,
32'b00000000111111111111000000000000,
32'b00000000111111111111000000000000,
32'b00000000111111111111000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b00001111111100000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111000000000000000000000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b11111111111111111111111100000000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00001111111111111111111100000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
         // code x07
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111111111111111111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b11111111000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000000000111111110000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000000001111111100000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000000011111111000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000111111110000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
        };

	assign data = ROM[addr];

endmodule  