module hexDriver (input  [3:0]  In0,
                  output logic [6:0]  Out0);
	
	always_comb
	begin
		unique case (In0)
	 	   4'b0000   : Out0 = 7'b0000001; // '0' b1000000 b0000001
	 	   4'b0001   : Out0 = 7'b1001111; // '1' b1111001 b1001111
		   4'b0010   : Out0 = 7'b0010010; // '2' b0100100 b0010010
	 	   4'b0011   : Out0 = 7'b0000110; // '3' b0110000 b0000110
	 	   4'b0100   : Out0 = 7'b1001100; // '4' b0011001 b1001100
		   4'b0101   : Out0 = 7'b0100100; // '5' b0010010 b0100100
	 	   4'b0110   : Out0 = 7'b0100000; // '6' b0000010 b0100000
	 	   4'b0111   : Out0 = 7'b0001111; // '7' b1111000 b0001111
	 	   4'b1000   : Out0 = 7'b0000000; // '8' b0000000 b0000000
		   4'b1001   : Out0 = 7'b0000100; // '9' b0010000 b0000100
	 	   4'b1010   : Out0 = 7'b0001000; // 'A' b0001000 b0001000
	 	   4'b1011   : Out0 = 7'b1100000; // 'b' b0000011 b1100000
	 	   4'b1100   : Out0 = 7'b0110001; // 'C' b1000110 b0110001
		   4'b1101   : Out0 = 7'b1000010; // 'd' b0100001 b1000010
	 	   4'b1110   : Out0 = 7'b0110000; // 'E' b0000110 b0110000
	 	   4'b1111   : Out0 = 7'b0111000; // 'F' b0001110 b0111000
	 	   default   : Out0 = 7'bX;
	  	 endcase
	end

endmodule